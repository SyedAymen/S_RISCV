module memory (
    input clk,
    output slow_clk
);
    assign slow_clk = clk;
endmodule
